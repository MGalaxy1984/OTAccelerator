module SenderTreeCluster
#(
  parameter TREE_NUM = 8,
  parameter AES_LATENCY
)
(
  input clk,
  input rst,
  input enable,
  input func,
  input [127:0] seed,
  input [127:0] delta,
  input [31:0] msg_index,
  output done,
  output reg [127:0] out
)

genvar i;
generate

endgenerate

endmodule