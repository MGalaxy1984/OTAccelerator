module BRAM_inst
#(parameter DATA_WIDTH=128,
  parameter ADDR_WIDTH=6)
(
  input [(DATA_WIDTH-1):0] data_in,
  input [(ADDR_WIDTH-1):0] read_addr, write_addr,
  input wr_en, clk,
  output logic [(DATA_WIDTH-1):0] data_out
);

(* ram_style = "block" *) reg [DATA_WIDTH-1:0] ram[2**ADDR_WIDTH-1:0];
// reg [ADDR_WIDTH-1:0] read_addr_reg;
   
always @ (posedge clk) begin
  // read_addr_reg <= read_addr; 
      
  if (wr_en) begin
    ram[write_addr] <= data_in;
  data_out <= ram[read_addr];
  end

end

// assign data_out = ram[read_addr_reg];
// assign data_out = ram[read_addr];

endmodule